module ysyx_25030077_IDU(
  input  [31:0] io_instruction,
  output [2:0]  io_imm_type,
  output [4:0]  io_rs1,
  output [4:0]  io_rs2,
  output [4:0]  io_rd,
  output [2:0]  io_data_control,
  output [3:0]  io_ALU_ctrl,
  output [3:0]  io_pc_next_type,
  output        is_break_out
);

  import "DPI-C" function bit is_break(input bit[31:0] instruction_in);
  assign is_break_out = is_break(io_instruction);

  wire [4:0] addi_Rs1 = io_instruction[19:15]; // @[module.scala 27:32]
  wire [4:0] addi_Rd = io_instruction[11:7]; // @[module.scala 28:32]
  wire [4:0] sltu_Rs2 = io_instruction[24:20]; // @[module.scala 75:33]
  wire [9:0] _isaddi_T_2 = {io_instruction[14:12],io_instruction[6:0]}; // @[Cat.scala 31:58]
  wire  isaddi = _isaddi_T_2 == 10'h13; // @[module.scala 256:64]
  wire  isxori = _isaddi_T_2 == 10'h213; // @[module.scala 257:64]
  wire  isori = _isaddi_T_2 == 10'h313; // @[module.scala 258:64]
  wire  isandi = _isaddi_T_2 == 10'h393; // @[module.scala 259:64]
  wire [15:0] _issrai_T_3 = {io_instruction[31:26],io_instruction[14:12],io_instruction[6:0]}; // @[Cat.scala 31:58]
  wire  issrai = _issrai_T_3 == 16'h4293; // @[module.scala 260:87]
  wire  issrli = _issrai_T_3 == 16'h293; // @[module.scala 261:87]
  wire  isslli = _issrai_T_3 == 16'h93; // @[module.scala 262:87]
  wire  issra = _issrai_T_3 == 16'h42b3; // @[module.scala 263:87]
  wire  issrl = _issrai_T_3 == 16'h2b3; // @[module.scala 264:87]
  wire  isbeq = _isaddi_T_2 == 10'h63; // @[module.scala 265:64]
  wire  isbne = _isaddi_T_2 == 10'he3; // @[module.scala 266:64]
  wire [16:0] _isadd_T_3 = {io_instruction[31:25],io_instruction[14:12],io_instruction[6:0]}; // @[Cat.scala 31:58]
  wire  isadd = _isadd_T_3 == 17'h33; // @[module.scala 267:87]
  wire  isxor = _isadd_T_3 == 17'h233; // @[module.scala 268:87]
  wire  isand = _isadd_T_3 == 17'h3b3; // @[module.scala 269:87]
  wire  isor = _isadd_T_3 == 17'h333; // @[module.scala 270:87]
  wire  issub = _isadd_T_3 == 17'h8033; // @[module.scala 271:87]
  wire  islui = io_instruction[6:0] == 7'h37; // @[module.scala 272:36]
  wire  isauipc = io_instruction[6:0] == 7'h17; // @[module.scala 273:38]
  wire  isjal = io_instruction[6:0] == 7'h6f; // @[module.scala 274:36]
  wire  isjalr = _isaddi_T_2 == 10'h67; // @[module.scala 275:65]
  wire  issw = _isaddi_T_2 == 10'h123; // @[module.scala 276:63]
  wire  isbge = _isaddi_T_2 == 10'h2e3; // @[module.scala 277:63]
  wire  isblt = _isaddi_T_2 == 10'h263; // @[module.scala 278:63]
  wire  isbltu = _isaddi_T_2 == 10'h363; // @[module.scala 279:63]
  wire  isbgeu = _isaddi_T_2 == 10'h3e3; // @[module.scala 280:63]
  wire  issb = _isaddi_T_2 == 10'h23; // @[module.scala 281:63]
  wire  issh = _isaddi_T_2 == 10'ha3; // @[module.scala 282:63]
  wire  islbu = _isaddi_T_2 == 10'h203; // @[module.scala 283:63]
  wire  islw = _isaddi_T_2 == 10'h103; // @[module.scala 284:63]
  wire  islh = _isaddi_T_2 == 10'h83; // @[module.scala 285:63]
  wire  islhu = _isaddi_T_2 == 10'h283; // @[module.scala 286:63]
  wire  issll = _isadd_T_3 == 17'hb3; // @[module.scala 287:86]
  wire  isslt = _isadd_T_3 == 17'h133; // @[module.scala 288:88]
  wire  issltu = _isadd_T_3 == 17'h1b3; // @[module.scala 289:88]
  wire  issltiu = _isaddi_T_2 == 10'h193; // @[module.scala 290:65]
  wire  isebreak = io_instruction == 32'h100073; // @[module.scala 291:34]
  wire [2:0] _io_imm_type_T = islbu ? 3'h1 : 3'h0; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_1 = islhu ? 3'h1 : _io_imm_type_T; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_2 = islh ? 3'h1 : _io_imm_type_T_1; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_3 = islw ? 3'h1 : _io_imm_type_T_2; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_4 = issh ? 3'h4 : _io_imm_type_T_3; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_5 = issb ? 3'h4 : _io_imm_type_T_4; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_6 = issw ? 3'h4 : _io_imm_type_T_5; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_7 = isjalr ? 3'h3 : _io_imm_type_T_6; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_8 = isjal ? 3'h3 : _io_imm_type_T_7; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_9 = isauipc ? 3'h2 : _io_imm_type_T_8; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_10 = islui ? 3'h2 : _io_imm_type_T_9; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_11 = issltiu ? 3'h1 : _io_imm_type_T_10; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_12 = isslli ? 3'h5 : _io_imm_type_T_11; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_13 = issrli ? 3'h5 : _io_imm_type_T_12; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_14 = issrai ? 3'h5 : _io_imm_type_T_13; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_15 = isandi ? 3'h1 : _io_imm_type_T_14; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_16 = isori ? 3'h1 : _io_imm_type_T_15; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_17 = isxori ? 3'h1 : _io_imm_type_T_16; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T = isslt ? addi_Rs1 : 5'h0; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_1 = issltu ? addi_Rs1 : _io_rs1_T; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_2 = isbne ? addi_Rs1 : _io_rs1_T_1; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_3 = isbgeu ? addi_Rs1 : _io_rs1_T_2; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_4 = isbltu ? addi_Rs1 : _io_rs1_T_3; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_5 = isblt ? addi_Rs1 : _io_rs1_T_4; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_6 = isbge ? addi_Rs1 : _io_rs1_T_5; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_7 = isbeq ? addi_Rs1 : _io_rs1_T_6; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_8 = issub ? addi_Rs1 : _io_rs1_T_7; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_9 = isor ? addi_Rs1 : _io_rs1_T_8; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_10 = isxor ? addi_Rs1 : _io_rs1_T_9; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_11 = issrl ? addi_Rs1 : _io_rs1_T_10; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_12 = issra ? addi_Rs1 : _io_rs1_T_11; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_13 = issll ? addi_Rs1 : _io_rs1_T_12; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_14 = isand ? addi_Rs1 : _io_rs1_T_13; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_15 = isadd ? addi_Rs1 : _io_rs1_T_14; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_16 = islbu ? addi_Rs1 : _io_rs1_T_15; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_17 = islhu ? addi_Rs1 : _io_rs1_T_16; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_18 = islh ? addi_Rs1 : _io_rs1_T_17; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_19 = islw ? addi_Rs1 : _io_rs1_T_18; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_20 = issh ? addi_Rs1 : _io_rs1_T_19; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_21 = issb ? addi_Rs1 : _io_rs1_T_20; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_22 = issw ? addi_Rs1 : _io_rs1_T_21; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_23 = isjalr ? addi_Rs1 : _io_rs1_T_22; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_24 = issltiu ? addi_Rs1 : _io_rs1_T_23; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_25 = isslli ? addi_Rs1 : _io_rs1_T_24; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_26 = issrli ? addi_Rs1 : _io_rs1_T_25; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_27 = issrai ? addi_Rs1 : _io_rs1_T_26; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_28 = isandi ? addi_Rs1 : _io_rs1_T_27; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_29 = isori ? addi_Rs1 : _io_rs1_T_28; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_30 = isxori ? addi_Rs1 : _io_rs1_T_29; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T = isslt ? sltu_Rs2 : 5'h0; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_1 = issltu ? sltu_Rs2 : _io_rs2_T; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_2 = isbne ? sltu_Rs2 : _io_rs2_T_1; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_3 = isbgeu ? sltu_Rs2 : _io_rs2_T_2; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_4 = isbltu ? sltu_Rs2 : _io_rs2_T_3; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_5 = isblt ? sltu_Rs2 : _io_rs2_T_4; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_6 = isbge ? sltu_Rs2 : _io_rs2_T_5; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_7 = isbeq ? sltu_Rs2 : _io_rs2_T_6; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_8 = issub ? sltu_Rs2 : _io_rs2_T_7; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_9 = isor ? sltu_Rs2 : _io_rs2_T_8; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_10 = isxor ? sltu_Rs2 : _io_rs2_T_9; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_11 = issrl ? sltu_Rs2 : _io_rs2_T_10; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_12 = issra ? sltu_Rs2 : _io_rs2_T_11; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_13 = issll ? sltu_Rs2 : _io_rs2_T_12; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_14 = isand ? sltu_Rs2 : _io_rs2_T_13; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_15 = isadd ? sltu_Rs2 : _io_rs2_T_14; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_16 = issh ? sltu_Rs2 : _io_rs2_T_15; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_17 = issb ? sltu_Rs2 : _io_rs2_T_16; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T = isslt ? addi_Rd : 5'h0; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_1 = issltu ? addi_Rd : _io_rd_T; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_2 = issub ? addi_Rd : _io_rd_T_1; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_3 = isor ? addi_Rd : _io_rd_T_2; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_4 = isxor ? addi_Rd : _io_rd_T_3; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_5 = issrl ? addi_Rd : _io_rd_T_4; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_6 = issra ? addi_Rd : _io_rd_T_5; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_7 = issll ? addi_Rd : _io_rd_T_6; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_8 = isand ? addi_Rd : _io_rd_T_7; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_9 = isadd ? addi_Rd : _io_rd_T_8; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_10 = islbu ? addi_Rd : _io_rd_T_9; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_11 = islhu ? addi_Rd : _io_rd_T_10; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_12 = islh ? addi_Rd : _io_rd_T_11; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_13 = islw ? addi_Rd : _io_rd_T_12; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_14 = isjalr ? addi_Rd : _io_rd_T_13; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_15 = isjal ? addi_Rd : _io_rd_T_14; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_16 = isauipc ? addi_Rd : _io_rd_T_15; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_17 = islui ? addi_Rd : _io_rd_T_16; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_18 = issltiu ? addi_Rd : _io_rd_T_17; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_19 = isslli ? addi_Rd : _io_rd_T_18; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_20 = issrli ? addi_Rd : _io_rd_T_19; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_21 = issrai ? addi_Rd : _io_rd_T_20; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_22 = isandi ? addi_Rd : _io_rd_T_21; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_23 = isori ? addi_Rd : _io_rd_T_22; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_24 = isxori ? addi_Rd : _io_rd_T_23; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T = issltu ? 5'h2 : 5'h0; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_1 = isslt ? 5'ha : _io_ALU_ctrl_T; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_2 = isbne ? 5'h0 : _io_ALU_ctrl_T_1; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_3 = isbgeu ? 5'h0 : _io_ALU_ctrl_T_2; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_4 = isbltu ? 5'h0 : _io_ALU_ctrl_T_3; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_5 = isblt ? 5'h0 : _io_ALU_ctrl_T_4; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_6 = isbge ? 5'h0 : _io_ALU_ctrl_T_5; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_7 = isbeq ? 5'h0 : _io_ALU_ctrl_T_6; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_8 = issub ? 5'h1 : _io_ALU_ctrl_T_7; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_9 = isor ? 5'h3 : _io_ALU_ctrl_T_8; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_10 = isxor ? 5'h4 : _io_ALU_ctrl_T_9; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_11 = issrl ? 5'h9 : _io_ALU_ctrl_T_10; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_12 = issra ? 5'h5 : _io_ALU_ctrl_T_11; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_13 = issll ? 5'h8 : _io_ALU_ctrl_T_12; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_14 = isand ? 5'h6 : _io_ALU_ctrl_T_13; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_15 = isadd ? 5'h0 : _io_ALU_ctrl_T_14; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_16 = islbu ? 5'h0 : _io_ALU_ctrl_T_15; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_17 = islhu ? 5'h0 : _io_ALU_ctrl_T_16; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_18 = islh ? 5'h0 : _io_ALU_ctrl_T_17; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_19 = islw ? 5'h0 : _io_ALU_ctrl_T_18; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_20 = issh ? 5'h0 : _io_ALU_ctrl_T_19; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_21 = issb ? 5'h0 : _io_ALU_ctrl_T_20; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_22 = issw ? 5'h0 : _io_ALU_ctrl_T_21; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_23 = isjalr ? 5'h0 : _io_ALU_ctrl_T_22; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_24 = isjal ? 5'h0 : _io_ALU_ctrl_T_23; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_25 = isauipc ? 5'h0 : _io_ALU_ctrl_T_24; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_26 = islui ? 5'h0 : _io_ALU_ctrl_T_25; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_27 = issltiu ? 5'h2 : _io_ALU_ctrl_T_26; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_28 = isslli ? 5'h8 : _io_ALU_ctrl_T_27; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_29 = issrli ? 5'h9 : _io_ALU_ctrl_T_28; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_30 = issrai ? 5'h5 : _io_ALU_ctrl_T_29; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_31 = isandi ? 5'h6 : _io_ALU_ctrl_T_30; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_32 = isori ? 5'h3 : _io_ALU_ctrl_T_31; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_33 = isxori ? 5'h4 : _io_ALU_ctrl_T_32; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_34 = isaddi ? 5'h0 : _io_ALU_ctrl_T_33; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T = issltu ? 3'h3 : 3'h0; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_1 = isslt ? 3'h3 : _io_data_control_T; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_2 = isbne ? 3'h0 : _io_data_control_T_1; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_3 = isbgeu ? 3'h0 : _io_data_control_T_2; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_4 = isbltu ? 3'h0 : _io_data_control_T_3; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_5 = isblt ? 3'h0 : _io_data_control_T_4; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_6 = isbge ? 3'h0 : _io_data_control_T_5; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_7 = isbeq ? 3'h0 : _io_data_control_T_6; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_8 = issub ? 3'h3 : _io_data_control_T_7; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_9 = isor ? 3'h3 : _io_data_control_T_8; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_10 = isxor ? 3'h3 : _io_data_control_T_9; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_11 = issrl ? 3'h3 : _io_data_control_T_10; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_12 = issra ? 3'h3 : _io_data_control_T_11; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_13 = issll ? 3'h3 : _io_data_control_T_12; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_14 = isand ? 3'h3 : _io_data_control_T_13; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_15 = isadd ? 3'h3 : _io_data_control_T_14; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_16 = islbu ? 3'h2 : _io_data_control_T_15; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_17 = islhu ? 3'h2 : _io_data_control_T_16; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_18 = islh ? 3'h2 : _io_data_control_T_17; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_19 = islw ? 3'h2 : _io_data_control_T_18; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_20 = issh ? 3'h0 : _io_data_control_T_19; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_21 = issb ? 3'h0 : _io_data_control_T_20; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_22 = issw ? 3'h0 : _io_data_control_T_21; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_23 = isjalr ? 3'h1 : _io_data_control_T_22; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_24 = isjal ? 3'h1 : _io_data_control_T_23; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T = issltiu ? 4'h0 : 4'h3; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_1 = isslt ? 4'h0 : _io_pc_next_type_T; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_2 = issltu ? 4'h0 : _io_pc_next_type_T_1; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_3 = isbne ? 4'h5 : _io_pc_next_type_T_2; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_4 = isbgeu ? 4'h8 : _io_pc_next_type_T_3; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_5 = isbltu ? 4'ha : _io_pc_next_type_T_4; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_6 = isblt ? 4'h9 : _io_pc_next_type_T_5; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_7 = isbge ? 4'h7 : _io_pc_next_type_T_6; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_8 = isbeq ? 4'h6 : _io_pc_next_type_T_7; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_9 = issub ? 4'h0 : _io_pc_next_type_T_8; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_10 = isor ? 4'h0 : _io_pc_next_type_T_9; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_11 = isxor ? 4'h0 : _io_pc_next_type_T_10; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_12 = issrl ? 4'h0 : _io_pc_next_type_T_11; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_13 = issra ? 4'h0 : _io_pc_next_type_T_12; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_14 = issll ? 4'h0 : _io_pc_next_type_T_13; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_15 = isand ? 4'h0 : _io_pc_next_type_T_14; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_16 = isadd ? 4'h0 : _io_pc_next_type_T_15; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_17 = islbu ? 4'h0 : _io_pc_next_type_T_16; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_18 = islhu ? 4'h0 : _io_pc_next_type_T_17; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_19 = islh ? 4'h0 : _io_pc_next_type_T_18; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_20 = islw ? 4'h0 : _io_pc_next_type_T_19; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_21 = isebreak ? 4'h4 : _io_pc_next_type_T_20; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_22 = issh ? 4'h0 : _io_pc_next_type_T_21; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_23 = issb ? 4'h0 : _io_pc_next_type_T_22; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_24 = issw ? 4'h0 : _io_pc_next_type_T_23; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_25 = isslli ? 4'h0 : _io_pc_next_type_T_24; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_26 = issrli ? 4'h0 : _io_pc_next_type_T_25; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_27 = issrai ? 4'h0 : _io_pc_next_type_T_26; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_28 = isandi ? 4'h0 : _io_pc_next_type_T_27; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_29 = isori ? 4'h0 : _io_pc_next_type_T_28; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_30 = isxori ? 4'h0 : _io_pc_next_type_T_29; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_31 = isaddi ? 4'h0 : _io_pc_next_type_T_30; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_32 = islui ? 4'h0 : _io_pc_next_type_T_31; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_33 = isauipc ? 4'h0 : _io_pc_next_type_T_32; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_34 = isjalr ? 4'h2 : _io_pc_next_type_T_33; // @[Mux.scala 101:16]
  assign io_imm_type = isaddi ? 3'h1 : _io_imm_type_T_17; // @[Mux.scala 101:16]
  assign io_rs1 = isaddi ? addi_Rs1 : _io_rs1_T_30; // @[Mux.scala 101:16]
  assign io_rs2 = issw ? sltu_Rs2 : _io_rs2_T_17; // @[Mux.scala 101:16]
  assign io_rd = isaddi ? addi_Rd : _io_rd_T_24; // @[Mux.scala 101:16]
  assign io_data_control = isauipc ? 3'h1 : _io_data_control_T_24; // @[Mux.scala 101:16]
  assign io_ALU_ctrl = _io_ALU_ctrl_T_34[3:0]; // @[module.scala 403:15]
  assign io_pc_next_type = isjal ? 4'h1 : _io_pc_next_type_T_34; // @[Mux.scala 101:16]
endmodule